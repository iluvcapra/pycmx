TITLE:   cdl_example02
FCM: NON-DROP FRAME 
000001  A205C016_220204_R24B             V     C        22:47:18:20 22:47:21:16 03:09:09:03 03:09:11:23 
*FROM CLIP NAME:  49D-3 
*ASC_SOP (0.98875 0.9878 0.98659)(-0.0008 0.00263 -0.00269)(0.9769 0.9767 0.97709) 
*ASC_SAT 1.0 
*SOURCE FILE: A205C016_220204_R24B 
000002  A238C007_220221_R24B             V     C        11:53:01:13 11:53:05:20 03:09:55:18 03:10:00:01 
*FROM CLIP NAME:  52B-7 
*ASC_SOP (1.05572 1.06914 1.05607)(-0.03004 -0.03044 -0.03044)(1.02112 1.01956 1.01707) 
*ASC_SAT 1.0 
*SOURCE FILE: A238C007_220221_R24B 
000004  A239C004_220221_R24B             V     C        15:19:53:22 15:19:55:02 03:10:00:01 03:10:01:05 
*FROM CLIP NAME:  52G-4* 
*ASC_SOP (1.00515 0.99542 0.9934)(-0.02412 -0.01467 -0.01351)(0.97348 0.97074 0.96887) 
*ASC_SAT 1.0 
*SOURCE FILE: A239C004_220221_R24B 
